library verilog;
use verilog.vl_types.all;
entity AES_top_vlg_vec_tst is
end AES_top_vlg_vec_tst;
