module GFM(A,B,C);

input [7:0] A,B;
output [7:0] C;

wire [7:0] w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13;

assign w0={8{A[7]}}&B;
assign w1={w0[6],w0[5],w0[4],w0[3],w0[2],w0[1],w0[0],1'b0}^{{8{w0[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w2=w1^{8{A[6]}}&B;
assign w3={w2[6],w2[5],w2[4],w2[3],w2[2],w2[1],w2[0],1'b0}^{{8{w2[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w4=w3^{8{A[5]}}&B;
assign w5={w4[6],w4[5],w4[4],w4[3],w4[2],w4[1],w4[0],1'b0}^{{8{w4[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w6=w5^{8{A[4]}}&B;
assign w7={w6[6],w6[5],w6[4],w6[3],w6[2],w6[1],w6[0],1'b0}^{{8{w6[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w8=w7^{8{A[3]}}&B;
assign w9={w8[6],w8[5],w8[4],w8[3],w8[2],w8[1],w8[0],1'b0}^{{8{w8[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w10=w9^{8{A[2]}}&B;
assign w11={w10[6],w10[5],w10[4],w10[3],w10[2],w10[1],w10[0],1'b0}^{{8{w10[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign w12=w11^{8{A[1]}}&B;
assign w13={w12[6],w12[5],w12[4],w12[3],w12[2],w12[1],w12[0],1'b0}^{{8{w12[7]}}&{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}};

assign C=w13^{8{A[0]}}&B;

endmodule
